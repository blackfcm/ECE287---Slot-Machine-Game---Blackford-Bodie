module character_rom(
    input  wire       clk,
    input  wire [7:0] ascii,   
    input  wire [3:0] row,     
    output reg  [7:0] pixels   
);

    
    reg [7:0] font[0:128*8-1];

    initial begin
        

        
        font[32*8+0]=8'b00000000;
        font[32*8+1]=8'b00000000;
        font[32*8+2]=8'b00000000;
        font[32*8+3]=8'b00000000;
        font[32*8+4]=8'b00000000;
        font[32*8+5]=8'b00000000;
        font[32*8+6]=8'b00000000;
        font[32*8+7]=8'b00000000;

        // F
        font["F"*8+0]=8'b11111110;
        font["F"*8+1]=8'b11111110;
        font["F"*8+2]=8'b11000000;
        font["F"*8+3]=8'b11000000;
        font["F"*8+4]=8'b11111100;
        font["F"*8+5]=8'b11111100;
        font["F"*8+6]=8'b11000000;
        font["F"*8+7]=8'b11000000;

        // o
        font["o"*8+0]=8'b00000000;
        font["o"*8+1]=8'b01111000;
        font["o"*8+2]=8'b11001100;
        font["o"*8+3]=8'b11001100;
        font["o"*8+4]=8'b11001100;
        font["o"*8+5]=8'b11001100;
        font["o"*8+6]=8'b01111000;
        font["o"*8+7]=8'b00000000;

        // r
        font["r"*8+0]=8'b00000000;
        font["r"*8+1]=8'b11111000;
        font["r"*8+2]=8'b11001100;
        font["r"*8+3]=8'b11000000;
        font["r"*8+4]=8'b11000000;
        font["r"*8+5]=8'b11000000;
        font["r"*8+6]=8'b11000000;
        font["r"*8+7]=8'b00000000;

        // t
        font["t"*8+0]=8'b00110000;
        font["t"*8+1]=8'b00110000;
        font["t"*8+2]=8'b11111100;
        font["t"*8+3]=8'b11111100;
        font["t"*8+4]=8'b00110000;
        font["t"*8+5]=8'b00110000;
        font["t"*8+6]=8'b00111100;
        font["t"*8+7]=8'b00000000;

        // u
        font["u"*8+0]=8'b00000000;
        font["u"*8+1]=8'b11001100;
        font["u"*8+2]=8'b11001100;
        font["u"*8+3]=8'b11001100;
        font["u"*8+4]=8'b11001100;
        font["u"*8+5]=8'b11001100;
        font["u"*8+6]=8'b01111100;
        font["u"*8+7]=8'b00000000;

        // n
        font["n"*8+0]=8'b00000000;
        font["n"*8+1]=8'b11111000;
        font["n"*8+2]=8'b11001100;
        font["n"*8+3]=8'b11001100;
        font["n"*8+4]=8'b11001100;
        font["n"*8+5]=8'b11001100;
        font["n"*8+6]=8'b11001100;
        font["n"*8+7]=8'b00000000;

        // e
        font["e"*8+0]=8'b00000000;
        font["e"*8+1]=8'b01111000;
        font["e"*8+2]=8'b11001100;
        font["e"*8+3]=8'b11111100;
        font["e"*8+4]=8'b11000000;
        font["e"*8+5]=8'b11000000;
        font["e"*8+6]=8'b01111100;
        font["e"*8+7]=8'b00000000;

        // z
        font["z"*8+0]=8'b00000000;
        font["z"*8+1]=8'b11111100;
        font["z"*8+2]=8'b00001100;
        font["z"*8+3]=8'b00111000;
        font["z"*8+4]=8'b01100000;
        font["z"*8+5]=8'b11000000;
        font["z"*8+6]=8'b11111100;
        font["z"*8+7]=8'b00000000;

        // y
        font["y"*8+0]=8'b00000000;
        font["y"*8+1]=8'b11001100;
        font["y"*8+2]=8'b11001100;
        font["y"*8+3]=8'b11001100;
        font["y"*8+4]=8'b01111100;
        font["y"*8+5]=8'b00001100;
        font["y"*8+6]=8'b11111000;
        font["y"*8+7]=8'b00000000;
		  
		  // Y
			font["Y"*8+0] = 8'b11000110;
			font["Y"*8+1] = 8'b11000110;
			font["Y"*8+2] = 8'b01101100;
			font["Y"*8+3] = 8'b00111000;
			font["Y"*8+4] = 8'b00111000;
			font["Y"*8+5] = 8'b00111000;
			font["Y"*8+6] = 8'b00111000;
			font["Y"*8+7] = 8'b00000000;
			
			// O
			font["O"*8+0] = 8'b00111000;
			font["O"*8+1] = 8'b01101100;
			font["O"*8+2] = 8'b11000110;
			font["O"*8+3] = 8'b11000110;
			font["O"*8+4] = 8'b11000110;
			font["O"*8+5] = 8'b11000110;
			font["O"*8+6] = 8'b01101100;
			font["O"*8+7] = 8'b00111000;
			
			// U
			font["U"*8+0] = 8'b11000110;
			font["U"*8+1] = 8'b11000110;
			font["U"*8+2] = 8'b11000110;
			font["U"*8+3] = 8'b11000110;
			font["U"*8+4] = 8'b11000110;
			font["U"*8+5] = 8'b11000110;
			font["U"*8+6] = 8'b01111100;
			font["U"*8+7] = 8'b00000000;
			
			// W
			font["W"*8+0] = 8'b11000110;
			font["W"*8+1] = 8'b11000110;
			font["W"*8+2] = 8'b11000110;
			font["W"*8+3] = 8'b11000110;
			font["W"*8+4] = 8'b11010110;
			font["W"*8+5] = 8'b11111110;
			font["W"*8+6] = 8'b01101100;
			font["W"*8+7] = 8'b00000000;

			// I
			font["I"*8+0] = 8'b11111110;
			font["I"*8+1] = 8'b00110000;
			font["I"*8+2] = 8'b00110000;
			font["I"*8+3] = 8'b00110000;
			font["I"*8+4] = 8'b00110000;
			font["I"*8+5] = 8'b00110000;
			font["I"*8+6] = 8'b11111110;
			font["I"*8+7] = 8'b00000000;
			
			// N
			font["N"*8+0] = 8'b11000110;
			font["N"*8+1] = 8'b11100110;
			font["N"*8+2] = 8'b11110110;
			font["N"*8+3] = 8'b11011110;
			font["N"*8+4] = 8'b11001110;
			font["N"*8+5] = 8'b11000110;
			font["N"*8+6] = 8'b11000110;
			font["N"*8+7] = 8'b00000000;
			
			// !
			font["!"*8+0] = 8'b00110000;
			font["!"*8+1] = 8'b00110000;
			font["!"*8+2] = 8'b00110000;
			font["!"*8+3] = 8'b00110000;
			font["!"*8+4] = 8'b00110000;
			font["!"*8+5] = 8'b00000000;
			font["!"*8+6] = 8'b00110000;
			font["!"*8+7] = 8'b00000000;

			// Letters for BET
			font["B"*8+0] = 8'b11111100;
			font["B"*8+1] = 8'b11000110;
			font["B"*8+2] = 8'b11000110;
			font["B"*8+3] = 8'b11111100;
			font["B"*8+4] = 8'b11000110;
			font["B"*8+5] = 8'b11000110;
			font["B"*8+6] = 8'b11111100;
			font["B"*8+7] = 8'b00000000;

			font["E"*8+0] = 8'b11111110;
			font["E"*8+1] = 8'b11000000;
			font["E"*8+2] = 8'b11000000;
			font["E"*8+3] = 8'b11111100;
			font["E"*8+4] = 8'b11000000;
			font["E"*8+5] = 8'b11000000;
			font["E"*8+6] = 8'b11111110;
			font["E"*8+7] = 8'b00000000;

			font["T"*8+0] = 8'b11111110;
			font["T"*8+1] = 8'b00110000;
			font["T"*8+2] = 8'b00110000;
			font["T"*8+3] = 8'b00110000;
			font["T"*8+4] = 8'b00110000;
			font["T"*8+5] = 8'b00110000;
			font["T"*8+6] = 8'b00110000;
			font["T"*8+7] = 8'b00000000;

			// Letters for PAYOUT
			font["P"*8+0] = 8'b11111100;
			font["P"*8+1] = 8'b11000110;
			font["P"*8+2] = 8'b11000110;
			font["P"*8+3] = 8'b11111100;
			font["P"*8+4] = 8'b11000000;
			font["P"*8+5] = 8'b11000000;
			font["P"*8+6] = 8'b11000000;
			font["P"*8+7] = 8'b00000000;

			font["A"*8+0] = 8'b01111100;
			font["A"*8+1] = 8'b11000110;
			font["A"*8+2] = 8'b11000110;
			font["A"*8+3] = 8'b11111110;
			font["A"*8+4] = 8'b11000110;
			font["A"*8+5] = 8'b11000110;
			font["A"*8+6] = 8'b11000110;
			font["A"*8+7] = 8'b00000000;

			font["Y"*8+0] = 8'b11000110;
			font["Y"*8+1] = 8'b11000110;
			font["Y"*8+2] = 8'b01101100;
			font["Y"*8+3] = 8'b00111000;
			font["Y"*8+4] = 8'b00111000;
			font["Y"*8+5] = 8'b00111000;
			font["Y"*8+6] = 8'b00111000;
			font["Y"*8+7] = 8'b00000000;

			font["O"*8+0] = 8'b00111000;
			font["O"*8+1] = 8'b01101100;
			font["O"*8+2] = 8'b11000110;
			font["O"*8+3] = 8'b11000110;
			font["O"*8+4] = 8'b11000110;
			font["O"*8+5] = 8'b11000110;
			font["O"*8+6] = 8'b01101100;
			font["O"*8+7] = 8'b00111000;

			font["U"*8+0] = 8'b11000110;
			font["U"*8+1] = 8'b11000110;
			font["U"*8+2] = 8'b11000110;
			font["U"*8+3] = 8'b11000110;
			font["U"*8+4] = 8'b11000110;
			font["U"*8+5] = 8'b11000110;
			font["U"*8+6] = 8'b01111100;
			font["U"*8+7] = 8'b00000000;

			// Digits 0-9
			font["0"*8+0] = 8'b01111100;
			font["0"*8+1] = 8'b11000110;
			font["0"*8+2] = 8'b11001110;
			font["0"*8+3] = 8'b11010110;
			font["0"*8+4] = 8'b11100110;
			font["0"*8+5] = 8'b11000110;
			font["0"*8+6] = 8'b01111100;
			font["0"*8+7] = 8'b00000000;

			font["1"*8+0] = 8'b00110000;
			font["1"*8+1] = 8'b01110000;
			font["1"*8+2] = 8'b00110000;
			font["1"*8+3] = 8'b00110000;
			font["1"*8+4] = 8'b00110000;
			font["1"*8+5] = 8'b00110000;
			font["1"*8+6] = 8'b11111100;
			font["1"*8+7] = 8'b00000000;
			
			font["2"*8+0] = 8'b01111100;
			font["2"*8+1] = 8'b11000110;
			font["2"*8+2] = 8'b00000110;
			font["2"*8+3] = 8'b00001100;
			font["2"*8+4] = 8'b00110000;
			font["2"*8+5] = 8'b01100000;
			font["2"*8+6] = 8'b11111110;
			font["2"*8+7] = 8'b00000000;
			
			font["3"*8+0] = 8'b01111100;
			font["3"*8+1] = 8'b11000110;
			font["3"*8+2] = 8'b00000110;
			font["3"*8+3] = 8'b00111100;
			font["3"*8+4] = 8'b00000110;
			font["3"*8+5] = 8'b11000110;
			font["3"*8+6] = 8'b01111100;
			font["3"*8+7] = 8'b00000000;
		
			font["4"*8+0] = 8'b00001100;
			font["4"*8+1] = 8'b00011100;
			font["4"*8+2] = 8'b00101100;
			font["4"*8+3] = 8'b01001100;
			font["4"*8+4] = 8'b11111110;
			font["4"*8+5] = 8'b00001100;
			font["4"*8+6] = 8'b00001100;
			font["4"*8+7] = 8'b00000000;
			
			font["5"*8+0] = 8'b11111110;
			font["5"*8+1] = 8'b11000000;
			font["5"*8+2] = 8'b11111100;
			font["5"*8+3] = 8'b00000110;
			font["5"*8+4] = 8'b00000110;
			font["5"*8+5] = 8'b11000110;
			font["5"*8+6] = 8'b01111100;
			font["5"*8+7] = 8'b00000000;
			
			font["6"*8+0] = 8'b01111100;
			font["6"*8+1] = 8'b11000110;
			font["6"*8+2] = 8'b11000000;
			font["6"*8+3] = 8'b11111100;
			font["6"*8+4] = 8'b11000110;
			font["6"*8+5] = 8'b11000110;
			font["6"*8+6] = 8'b01111100;
			font["6"*8+7] = 8'b00000000;
			
			font["7"*8+0] = 8'b11111110;
			font["7"*8+1] = 8'b00000110;
			font["7"*8+2] = 8'b00001100;
			font["7"*8+3] = 8'b00011000;
			font["7"*8+4] = 8'b00110000;
			font["7"*8+5] = 8'b01100000;
			font["7"*8+6] = 8'b01100000;
			font["7"*8+7] = 8'b00000000;
			
			font["8"*8+0] = 8'b01111100;
			font["8"*8+1] = 8'b11000110;
			font["8"*8+2] = 8'b11000110;
			font["8"*8+3] = 8'b01111100;
			font["8"*8+4] = 8'b11000110;
			font["8"*8+5] = 8'b11000110;
			font["8"*8+6] = 8'b01111100;
			font["8"*8+7] = 8'b00000000;

		font["9"*8+0] = 8'b01111100;
		font["9"*8+1] = 8'b11000110;
		font["9"*8+2] = 8'b11000110;
		font["9"*8+3] = 8'b01111110;
		font["9"*8+4] = 8'b00000110;
		font["9"*8+5] = 8'b11000110;
		font["9"*8+6] = 8'b01111100;
		font["9"*8+7] = 8'b00000000;
    end

    always @(posedge clk)
        pixels <= font[ascii*8 + row];

endmodule
